// tb meant to ensure connection between caches work
module l1d_llc_tb (
    // Input signals
    input logic clk,
    input logic rst_N,

    // L1D cache interface inputs
    
    // L1D cache interface outputs

);


endmodule
