// adjust refresh param based on the actual clock, currently assuming 1 GHz clock => 64 ms = 64,000,000 ns
module refresh_timer #(
    parameter int REFRESH = 64_000_000
) (
    input logic clk_in,
    input logic rst_in,
    output logic refresh
);
    localparam WIDTH = $clog2(REFRESH)
    logic [WIDTH-1:0] count;
    always_ff @(posedge clk or posedge rst_in) begin
        if (rst_in) begin
            count <= 0;
            refresh <= 0;
        end else if (count == REFRESH - 1) begin
            count <= 0;
            refresh <= ~refresh;
        end else begin
            count <= count + 1;
        end
    end 
endmodule : refresh_timer

module auto_refresh #(
    parameter int BANK_GROUPS = 2,
    parameter int BANKS_PER_GROUP = 4,       // banks per group
    parameter int ROW_BITS = 8,    // bits to address rows
    parameter int ACTIVATION_LATENCY = 8,
    parameter int PRECHARGE_LATENCY = 5, 
    parameter int REFRESH_LATENCY = ACTIVATION_LATENCY + PRECHARGE_LATENCY,
    parameter int BANKS = BANK_GROUPS * BANKS_PER_GROUP
) (
    input logic clk_in,
    input logic rst_in,
    input logic valid_in, // if not valid ignore,
    output logic [$clog2(BANK_GROUPS)-1:0] bank_group_out,
    output logic [$clog2(BANKS_PER_GROUP)-1:0] bank_out,
    output logic [ROW_BITS-1:0] row_out,
    output logic valid_out
);
    // iterate through all banks then all rows
    localparam BANK_BITS = $clog2(BANKS_PER_GROUP);
    localparam BANK_GRP_BITS = $clog2(BANK_GROUPS);
    logic [ROW_BITS:0] _state;
    logic [3:0] state; // might need to parameterize this later
    always_ff @(posedge clk_in or posedge rst_in) begin
        if (rst_in) begin
            _state <= 0;
            state <= 0;
        end else begin
            if (state == 12) begin
                if (_state == 1 << ROW_BITS - 1) begin
                    _state <= 0;
                end else begin
                    _state <= _state + 1;
                end
                state <= 0;
            end else begin
                state <= state + 1;
            end
        end
    end

    always_comb begin
        valid_out = '0;
        row_out = '0;
        bank_out = '0;
        bank_group_out = '0;
        if (valid_in) begin
            if (state < $clog2(BANKS)) begin
                valid_out = 1'b1;
                row_out = _state;
                bank_out = state & {{{13-BANK_BITS}{1'b0}}, {BANK_BITS{1'b1}}};
                bank_group_out = (state >> BANK_BITS) & {{{13-BANK_GRP_BITS}{1'b0}}, {BANK_GRP_BITS{1'b1}}};
            end
        end
    end
endmodule: auto_refresh